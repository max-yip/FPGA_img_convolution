module color_filter (
	input	 logic			 clk,
	input  logic 		 	 rst,
	input  logic [11:0] 	 pixel_in,
	input  logic 		 	 in_ready,
	input  logic 		 	 veml_ready,
	input  logic [15:0] 	 parcel_colour, // to be defined
	output logic [11:0] 	 pixel_out,
	output logic 			 out_ready
);

	

endmodule