module vga_scaler (
	input  logic [11:0] data_in,
	input  logic pclk,
	input  logic ready, 
	input  logic rst,
	output logic [11:0] data_out
);










endmodule